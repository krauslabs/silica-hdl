module and_gate (a, b, y);
    input a;
    input b;
    output y;
    assign y = a & b;
endmodule